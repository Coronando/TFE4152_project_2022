*NAND Gate subcircuit


*subcurcuit nand gate
.subckt nand input_a input_b out

Vdd v_main gnd DC 1.0V

*PMOS params
.param L_pmos = 100n
.param W_pmos = 100n
*NMOS params
.param L_nmos = 100n
.param W_nmos = 100n

*Upper part of circuit defined
XM_Apmos v_main input_a v_out v_main pmos1v L=L_pmos W=W_pmos
XM_Bpmos v_main input_b v_out v_main pmos1v L=L_pmos W=W_pmos

*Lower part of circuit defined
XM_Anmos v_out input_a gnd gnd nmos1v L=L_nmos W=W_nmos
XM_Bnmos v_out input_b gnd gnd nmos1v L=L_nmos W=W_nmos

.ends nand