*3 input AND Gate by Sindre Nordtveit and Mathias Bj�nnes

*NB: For this file to work, it has to be included AFTER the NOT and NAND

.subckt and_pg_gate input_a input_b sel output v_main gnd

Xpg_pmos    v_main      sel         top         v_main  pmos1v L=L_pmos W=W_pmos

*Upper part of NAND circuit
XM_Apmos    top         input_a     and_out     top     pmos1v L=L_pmos W=W_pmos
XM_Bpmos    top         input_b     and_out     top     pmos1v L=L_pmos W=W_pmos
*Lower part of NAND defined
XM_Anmos    and_out     input_a     a_source    bottom     nmos1v L=L_nmos W=W_nmos
XM_Bnmos    a_source    input_b     bottom      bottom     nmos1v L=L_nmos W=W_nmos

*Inverter
Xinv_pmos   top         and_out     output      top        pmos1v L=L_pmos W=W_pmos
Xinv_nmos   output      and_out     bottom      bottom     nmos1v L=L_nmos W=W_nmos

Xpg_nmos    bottom      sel         gnd         gnd     nmos1v L=L_nmos W=W_nmos

.ends and_pg_gate