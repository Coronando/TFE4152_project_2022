module test(input logic hello, output logic bye);
endmodule